ENTITY Decoder IS
	PORT (
		INPUT : IN BIT_VECTOR(3 DOWNTO 0);
		OUTPUT : OUT BIT_VECTOR(6 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE Decoder_Arch OF Decoder IS
	SIGNAL NINPUT : BIT_VECTOR(3 DOWNTO 0);

BEGIN
	NINPUT(0) <= NOT INPUT(0);
	NINPUT(1) <= NOT INPUT(1);
	NINPUT(2) <= NOT INPUT(2);
	NINPUT(3) <= NOT INPUT(3);

	OUTPUT(0) <= (INPUT(0) OR INPUT(1) OR INPUT(2) OR NINPUT(3)) AND (INPUT(0) OR NINPUT(1) OR INPUT(2) OR INPUT(3));
	OUTPUT(1) <= (INPUT(0) OR NINPUT(1) OR INPUT(2) OR NINPUT(3)) AND (INPUT(0) OR NINPUT(1) OR NINPUT(2) OR INPUT(3));
	OUTPUT(2) <= INPUT(0) OR INPUT(1) OR NINPUT(2) OR INPUT(3);
	OUTPUT(3) <= (INPUT(0) OR INPUT(1) OR INPUT(2) OR NINPUT(3)) AND (INPUT(0) OR NINPUT(1) OR INPUT(2) OR INPUT(3)) AND (INPUT(0) OR NINPUT(1) OR NINPUT(2) OR NINPUT(3));
	OUTPUT(4) <= INPUT(1) AND INPUT(3);
	OUTPUT(5) <= (INPUT(0) OR INPUT(1) OR NINPUT(3)) AND (INPUT(0) OR NINPUT(2) OR NINPUT(3)) AND (INPUT(0) OR INPUT(1) OR NINPUT(2) OR INPUT(3));
	OUTPUT(6) <= (INPUT(0) OR INPUT(1) OR INPUT(2)) AND (INPUT(0) OR NINPUT(1) OR NINPUT(2) OR NINPUT(3));
	
END ARCHITECTURE;
